module reg (d, q, ena, clk);
				
input	reg ena, clk, d7, d6, d5, d4, d3, d2, d1, d0;
output wire 		  q7, q6, q5, q4, q3, q2, q1, q0;














endmodule				